// Copyright 2025 Google LLC
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

//----------------------------------------------------------------------------
// Description:covergroup for RV32M instruction
//----------------------------------------------------------------------------
covergroup cvgrp_RV32_M;

    	option.per_instance = 1;
        // base cover
	mul: coverpoint rv32m_trans.inst_name iff(rv32m_trans.trap==0) {
		bins b0 = {MUL};
		option.weight = 1;
	 }

	mulh: coverpoint rv32m_trans.inst_name iff(rv32m_trans.trap==0) {
		bins b0 = {MULH};
		option.weight = 1;
	 }

	mulhsu: coverpoint rv32m_trans.inst_name iff(rv32m_trans.trap==0) {
		bins b0 = {MULHSU};
		option.weight = 1;
	 }

	mulhu: coverpoint rv32m_trans.inst_name iff(rv32m_trans.trap==0) {
		bins b0 = {MULHU};
		option.weight = 1;
	 }

	div: coverpoint rv32m_trans.inst_name iff(rv32m_trans.trap==0) {
		bins b0 = {DIV};
		option.weight = 1;
	 }

	divu: coverpoint rv32m_trans.inst_name iff(rv32m_trans.trap==0) {
		bins b0 = {DIVU};
		option.weight = 1;
	 }

	rem: coverpoint rv32m_trans.inst_name iff(rv32m_trans.trap==0) {
		bins b0 = {REM};
		option.weight = 1;
	 }

	remu: coverpoint rv32m_trans.inst_name iff(rv32m_trans.trap==0) {
		bins b0 = {REMU};
		option.weight = 1;
	 }

	//RD (GPR) register assignment,x0 always 0
	rd_addr: coverpoint rv32m_trans.rd_addr iff(rv32m_trans.trap==0) {
		bins b0 = {0};
		bins b1 = {1};
		bins b2 = {2};
		bins b3 = {3};
		bins b4 = {4};
		bins b5 = {5};
		bins b6 = {6};
		bins b7 = {7};
		bins b8 = {8};
		bins b9 = {9};
		bins b10 = {10};
		bins b11 = {11};
		bins b12 = {12};
		bins b13 = {13};
		bins b14 = {14};
		bins b15 = {15};
		bins b16 = {16};
		bins b17 = {17};
		bins b18 = {18};
		bins b19 = {19};
		bins b20 = {20};
		bins b21 = {21};
		bins b22 = {22};
		bins b23 = {23};
		bins b24 = {24};
		bins b25 = {25};
		bins b26 = {26};
		bins b27 = {27};
		bins b28 = {28};
		bins b29 = {29};
		bins b30 = {30};
		bins b31 = {31};
		option.weight = 1;
	 }

	//RS1 (GPR) register assignment
	rs1_addr: coverpoint rv32m_trans.rs1_addr iff(rv32m_trans.trap==0) {
		bins b0 = {0};
		bins b1 = {1};
		bins b2 = {2};
		bins b3 = {3};
		bins b4 = {4};
		bins b5 = {5};
		bins b6 = {6};
		bins b7 = {7};
		bins b8 = {8};
		bins b9 = {9};
		bins b10 = {10};
		bins b11 = {11};
		bins b12 = {12};
		bins b13 = {13};
		bins b14 = {14};
		bins b15 = {15};
		bins b16 = {16};
		bins b17 = {17};
		bins b18 = {18};
		bins b19 = {19};
		bins b20 = {20};
		bins b21 = {21};
		bins b22 = {22};
		bins b23 = {23};
		bins b24 = {24};
		bins b25 = {25};
		bins b26 = {26};
		bins b27 = {27};
		bins b28 = {28};
		bins b29 = {29};
		bins b30 = {30};
		bins b31 = {31};
		option.weight = 1;
	 }

	//RS2 (GPR) register assignment
	rs2_addr: coverpoint rv32m_trans.rs2_addr iff(rv32m_trans.trap==0) {
		bins b0 = {0};
		bins b1 = {1};
		bins b2 = {2};
		bins b3 = {3};
		bins b4 = {4};
		bins b5 = {5};
		bins b6 = {6};
		bins b7 = {7};
		bins b8 = {8};
		bins b9 = {9};
		bins b10 = {10};
		bins b11 = {11};
		bins b12 = {12};
		bins b13 = {13};
		bins b14 = {14};
		bins b15 = {15};
		bins b16 = {16};
		bins b17 = {17};
		bins b18 = {18};
		bins b19 = {19};
		bins b20 = {20};
		bins b21 = {21};
		bins b22 = {22};
		bins b23 = {23};
		bins b24 = {24};
		bins b25 = {25};
		bins b26 = {26};
		bins b27 = {27};
		bins b28 = {28};
		bins b29 = {29};
		bins b30 = {30};
		bins b31 = {31};
		option.weight = 1;
	 }

	//RD toggle bits
	rd_val: coverpoint unsigned'(rv32m_trans.rd_val) iff(rv32m_trans.trap==0) {
		wildcard bins b_1_0_0 	= (32'b???????????????????????????????1=>32'b???????????????????????????????0);
		wildcard bins b_1_0_1 	= (32'b??????????????????????????????1?=>32'b??????????????????????????????0?);
		wildcard bins b_1_0_2 	= (32'b?????????????????????????????1??=>32'b?????????????????????????????0??);
		wildcard bins b_1_0_3 	= (32'b????????????????????????????1???=>32'b????????????????????????????0???);
		wildcard bins b_1_0_4 	= (32'b???????????????????????????1????=>32'b???????????????????????????0????);
		wildcard bins b_1_0_5 	= (32'b??????????????????????????1?????=>32'b??????????????????????????0?????);
		wildcard bins b_1_0_6 	= (32'b?????????????????????????1??????=>32'b?????????????????????????0??????);
		wildcard bins b_1_0_7 	= (32'b????????????????????????1???????=>32'b????????????????????????0???????);
		wildcard bins b_1_0_8 	= (32'b???????????????????????1????????=>32'b???????????????????????0????????);
		wildcard bins b_1_0_9 	= (32'b??????????????????????1?????????=>32'b??????????????????????0?????????);
		wildcard bins b_1_0_10 	= (32'b?????????????????????1??????????=>32'b?????????????????????0??????????);
		wildcard bins b_1_0_11 	= (32'b????????????????????1???????????=>32'b????????????????????0???????????);
		wildcard bins b_1_0_12 	= (32'b???????????????????1????????????=>32'b???????????????????0????????????);
		wildcard bins b_1_0_13 	= (32'b??????????????????1?????????????=>32'b??????????????????0?????????????);
		wildcard bins b_1_0_14 	= (32'b?????????????????1??????????????=>32'b?????????????????0??????????????);
		wildcard bins b_1_0_15 	= (32'b????????????????1???????????????=>32'b????????????????0???????????????);
		wildcard bins b_1_0_16 	= (32'b???????????????1????????????????=>32'b???????????????0????????????????);
		wildcard bins b_1_0_17 	= (32'b??????????????1?????????????????=>32'b??????????????0?????????????????);
		wildcard bins b_1_0_18 	= (32'b?????????????1??????????????????=>32'b?????????????0??????????????????);
		wildcard bins b_1_0_19 	= (32'b????????????1???????????????????=>32'b????????????0???????????????????);
		wildcard bins b_1_0_20 	= (32'b???????????1????????????????????=>32'b???????????0????????????????????);
		wildcard bins b_1_0_21 	= (32'b??????????1?????????????????????=>32'b??????????0?????????????????????);
		wildcard bins b_1_0_22 	= (32'b?????????1??????????????????????=>32'b?????????0??????????????????????);
		wildcard bins b_1_0_23 	= (32'b????????1???????????????????????=>32'b????????0???????????????????????);
		wildcard bins b_1_0_24 	= (32'b???????1????????????????????????=>32'b???????0????????????????????????);
		wildcard bins b_1_0_25 	= (32'b??????1?????????????????????????=>32'b??????0?????????????????????????);
		wildcard bins b_1_0_26 	= (32'b?????1??????????????????????????=>32'b?????0??????????????????????????);
		wildcard bins b_1_0_27 	= (32'b????1???????????????????????????=>32'b????0???????????????????????????);
		wildcard bins b_1_0_28 	= (32'b???1????????????????????????????=>32'b???0????????????????????????????);
		wildcard bins b_1_0_29 	= (32'b??1?????????????????????????????=>32'b??0?????????????????????????????);
		wildcard bins b_1_0_30 	= (32'b?1??????????????????????????????=>32'b?0??????????????????????????????);
		wildcard bins b_1_0_31 	= (32'b1???????????????????????????????=>32'b0???????????????????????????????);
		wildcard bins b_0_1_0 	= (32'b???????????????????????????????0=>32'b???????????????????????????????1);
		wildcard bins b_0_1_1 	= (32'b??????????????????????????????0?=>32'b??????????????????????????????1?);
		wildcard bins b_0_1_2 	= (32'b?????????????????????????????0??=>32'b?????????????????????????????1??);
		wildcard bins b_0_1_3 	= (32'b????????????????????????????0???=>32'b????????????????????????????1???);
		wildcard bins b_0_1_4 	= (32'b???????????????????????????0????=>32'b???????????????????????????1????);
		wildcard bins b_0_1_5 	= (32'b??????????????????????????0?????=>32'b??????????????????????????1?????);
		wildcard bins b_0_1_6 	= (32'b?????????????????????????0??????=>32'b?????????????????????????1??????);
		wildcard bins b_0_1_7 	= (32'b????????????????????????0???????=>32'b????????????????????????1???????);
		wildcard bins b_0_1_8 	= (32'b???????????????????????0????????=>32'b???????????????????????1????????);
		wildcard bins b_0_1_9 	= (32'b??????????????????????0?????????=>32'b??????????????????????1?????????);
		wildcard bins b_0_1_10 	= (32'b?????????????????????0??????????=>32'b?????????????????????1??????????);
		wildcard bins b_0_1_11 	= (32'b????????????????????0???????????=>32'b????????????????????1???????????);
		wildcard bins b_0_1_12 	= (32'b???????????????????0????????????=>32'b???????????????????1????????????);
		wildcard bins b_0_1_13 	= (32'b??????????????????0?????????????=>32'b??????????????????1?????????????);
		wildcard bins b_0_1_14 	= (32'b?????????????????0??????????????=>32'b?????????????????1??????????????);
		wildcard bins b_0_1_15 	= (32'b????????????????0???????????????=>32'b????????????????1???????????????);
		wildcard bins b_0_1_16 	= (32'b???????????????0????????????????=>32'b???????????????1????????????????);
		wildcard bins b_0_1_17 	= (32'b??????????????0?????????????????=>32'b??????????????1?????????????????);
		wildcard bins b_0_1_18 	= (32'b?????????????0??????????????????=>32'b?????????????1??????????????????);
		wildcard bins b_0_1_19 	= (32'b????????????0???????????????????=>32'b????????????1???????????????????);
		wildcard bins b_0_1_20 	= (32'b???????????0????????????????????=>32'b???????????1????????????????????);
		wildcard bins b_0_1_21 	= (32'b??????????0?????????????????????=>32'b??????????1?????????????????????);
		wildcard bins b_0_1_22 	= (32'b?????????0??????????????????????=>32'b?????????1??????????????????????);
		wildcard bins b_0_1_23 	= (32'b????????0???????????????????????=>32'b????????1???????????????????????);
		wildcard bins b_0_1_24 	= (32'b???????0????????????????????????=>32'b???????1????????????????????????);
		wildcard bins b_0_1_25 	= (32'b??????0?????????????????????????=>32'b??????1?????????????????????????);
		wildcard bins b_0_1_26 	= (32'b?????0??????????????????????????=>32'b?????1??????????????????????????);
		wildcard bins b_0_1_27 	= (32'b????0???????????????????????????=>32'b????1???????????????????????????);
		wildcard bins b_0_1_28 	= (32'b???0????????????????????????????=>32'b???1????????????????????????????);
		wildcard bins b_0_1_29 	= (32'b??0?????????????????????????????=>32'b??1?????????????????????????????);
		wildcard bins b_0_1_30 	= (32'b?0??????????????????????????????=>32'b?1??????????????????????????????);
		wildcard bins b_0_1_31 	= (32'b0???????????????????????????????=>32'b1???????????????????????????????);
		option.weight = 1;
	 }

	//RD special values
	rd_sp_val: coverpoint unsigned'(rv32m_trans.rd_val) iff(rv32m_trans.trap==0) {
		bins b0 = {32'b0};
		bins b1 = {32'b00000000000000000000000000000001};
		bins b2 = {32'b11111111111111111111111111111111};
		bins b3 = {32'b01111111111111111111111111111111};
		bins b4 = {32'b10000000000000000000000000000000};
		bins b5 = {32'b10000000000000000000000000000001};
		option.weight = 1;
	 }

	//RD value sign
	rd_val_sign: coverpoint rv32m_trans.rd_val iff(rv32m_trans.trap==0) {
		bins b0 = {[$:-1]};
		bins b1 = {[1:$]};
		option.weight = 1;
	 }

	//RS1 toggle bits
	rs1_val: coverpoint unsigned'(rv32m_trans.rs1_val) iff(rv32m_trans.trap==0) {
		wildcard bins b_1_0_0 	= (32'b???????????????????????????????1=>32'b???????????????????????????????0);
		wildcard bins b_1_0_1 	= (32'b??????????????????????????????1?=>32'b??????????????????????????????0?);
		wildcard bins b_1_0_2 	= (32'b?????????????????????????????1??=>32'b?????????????????????????????0??);
		wildcard bins b_1_0_3 	= (32'b????????????????????????????1???=>32'b????????????????????????????0???);
		wildcard bins b_1_0_4 	= (32'b???????????????????????????1????=>32'b???????????????????????????0????);
		wildcard bins b_1_0_5 	= (32'b??????????????????????????1?????=>32'b??????????????????????????0?????);
		wildcard bins b_1_0_6 	= (32'b?????????????????????????1??????=>32'b?????????????????????????0??????);
		wildcard bins b_1_0_7 	= (32'b????????????????????????1???????=>32'b????????????????????????0???????);
		wildcard bins b_1_0_8 	= (32'b???????????????????????1????????=>32'b???????????????????????0????????);
		wildcard bins b_1_0_9 	= (32'b??????????????????????1?????????=>32'b??????????????????????0?????????);
		wildcard bins b_1_0_10 	= (32'b?????????????????????1??????????=>32'b?????????????????????0??????????);
		wildcard bins b_1_0_11 	= (32'b????????????????????1???????????=>32'b????????????????????0???????????);
		wildcard bins b_1_0_12 	= (32'b???????????????????1????????????=>32'b???????????????????0????????????);
		wildcard bins b_1_0_13 	= (32'b??????????????????1?????????????=>32'b??????????????????0?????????????);
		wildcard bins b_1_0_14 	= (32'b?????????????????1??????????????=>32'b?????????????????0??????????????);
		wildcard bins b_1_0_15 	= (32'b????????????????1???????????????=>32'b????????????????0???????????????);
		wildcard bins b_1_0_16 	= (32'b???????????????1????????????????=>32'b???????????????0????????????????);
		wildcard bins b_1_0_17 	= (32'b??????????????1?????????????????=>32'b??????????????0?????????????????);
		wildcard bins b_1_0_18 	= (32'b?????????????1??????????????????=>32'b?????????????0??????????????????);
		wildcard bins b_1_0_19 	= (32'b????????????1???????????????????=>32'b????????????0???????????????????);
		wildcard bins b_1_0_20 	= (32'b???????????1????????????????????=>32'b???????????0????????????????????);
		wildcard bins b_1_0_21 	= (32'b??????????1?????????????????????=>32'b??????????0?????????????????????);
		wildcard bins b_1_0_22 	= (32'b?????????1??????????????????????=>32'b?????????0??????????????????????);
		wildcard bins b_1_0_23 	= (32'b????????1???????????????????????=>32'b????????0???????????????????????);
		wildcard bins b_1_0_24 	= (32'b???????1????????????????????????=>32'b???????0????????????????????????);
		wildcard bins b_1_0_25 	= (32'b??????1?????????????????????????=>32'b??????0?????????????????????????);
		wildcard bins b_1_0_26 	= (32'b?????1??????????????????????????=>32'b?????0??????????????????????????);
		wildcard bins b_1_0_27 	= (32'b????1???????????????????????????=>32'b????0???????????????????????????);
		wildcard bins b_1_0_28 	= (32'b???1????????????????????????????=>32'b???0????????????????????????????);
		wildcard bins b_1_0_29 	= (32'b??1?????????????????????????????=>32'b??0?????????????????????????????);
		wildcard bins b_1_0_30 	= (32'b?1??????????????????????????????=>32'b?0??????????????????????????????);
		wildcard bins b_1_0_31 	= (32'b1???????????????????????????????=>32'b0???????????????????????????????);
		wildcard bins b_0_1_0 	= (32'b???????????????????????????????0=>32'b???????????????????????????????1);
		wildcard bins b_0_1_1 	= (32'b??????????????????????????????0?=>32'b??????????????????????????????1?);
		wildcard bins b_0_1_2 	= (32'b?????????????????????????????0??=>32'b?????????????????????????????1??);
		wildcard bins b_0_1_3 	= (32'b????????????????????????????0???=>32'b????????????????????????????1???);
		wildcard bins b_0_1_4 	= (32'b???????????????????????????0????=>32'b???????????????????????????1????);
		wildcard bins b_0_1_5 	= (32'b??????????????????????????0?????=>32'b??????????????????????????1?????);
		wildcard bins b_0_1_6 	= (32'b?????????????????????????0??????=>32'b?????????????????????????1??????);
		wildcard bins b_0_1_7 	= (32'b????????????????????????0???????=>32'b????????????????????????1???????);
		wildcard bins b_0_1_8 	= (32'b???????????????????????0????????=>32'b???????????????????????1????????);
		wildcard bins b_0_1_9 	= (32'b??????????????????????0?????????=>32'b??????????????????????1?????????);
		wildcard bins b_0_1_10 	= (32'b?????????????????????0??????????=>32'b?????????????????????1??????????);
		wildcard bins b_0_1_11 	= (32'b????????????????????0???????????=>32'b????????????????????1???????????);
		wildcard bins b_0_1_12 	= (32'b???????????????????0????????????=>32'b???????????????????1????????????);
		wildcard bins b_0_1_13 	= (32'b??????????????????0?????????????=>32'b??????????????????1?????????????);
		wildcard bins b_0_1_14 	= (32'b?????????????????0??????????????=>32'b?????????????????1??????????????);
		wildcard bins b_0_1_15 	= (32'b????????????????0???????????????=>32'b????????????????1???????????????);
		wildcard bins b_0_1_16 	= (32'b???????????????0????????????????=>32'b???????????????1????????????????);
		wildcard bins b_0_1_17 	= (32'b??????????????0?????????????????=>32'b??????????????1?????????????????);
		wildcard bins b_0_1_18 	= (32'b?????????????0??????????????????=>32'b?????????????1??????????????????);
		wildcard bins b_0_1_19 	= (32'b????????????0???????????????????=>32'b????????????1???????????????????);
		wildcard bins b_0_1_20 	= (32'b???????????0????????????????????=>32'b???????????1????????????????????);
		wildcard bins b_0_1_21 	= (32'b??????????0?????????????????????=>32'b??????????1?????????????????????);
		wildcard bins b_0_1_22 	= (32'b?????????0??????????????????????=>32'b?????????1??????????????????????);
		wildcard bins b_0_1_23 	= (32'b????????0???????????????????????=>32'b????????1???????????????????????);
		wildcard bins b_0_1_24 	= (32'b???????0????????????????????????=>32'b???????1????????????????????????);
		wildcard bins b_0_1_25 	= (32'b??????0?????????????????????????=>32'b??????1?????????????????????????);
		wildcard bins b_0_1_26 	= (32'b?????0??????????????????????????=>32'b?????1??????????????????????????);
		wildcard bins b_0_1_27 	= (32'b????0???????????????????????????=>32'b????1???????????????????????????);
		wildcard bins b_0_1_28 	= (32'b???0????????????????????????????=>32'b???1????????????????????????????);
		wildcard bins b_0_1_29 	= (32'b??0?????????????????????????????=>32'b??1?????????????????????????????);
		wildcard bins b_0_1_30 	= (32'b?0??????????????????????????????=>32'b?1??????????????????????????????);
		wildcard bins b_0_1_31 	= (32'b0???????????????????????????????=>32'b1???????????????????????????????);
		option.weight = 1;
	 }

	//RS1 special values
	rs1_sp_val: coverpoint unsigned'(rv32m_trans.rs1_val) iff(rv32m_trans.trap==0) {
		bins b0 = {32'b0};
		bins b1 = {32'b00000000000000000000000000000001};
		bins b2 = {32'b11111111111111111111111111111111};
		bins b3 = {32'b01111111111111111111111111111111};
		bins b4 = {32'b10000000000000000000000000000000};
		bins b5 = {32'b10000000000000000000000000000001};
		option.weight = 1;
	 }

	//RS1 value sign
	rs1_val_sign: coverpoint rv32m_trans.rs1_val iff(rv32m_trans.trap==0) {
		bins b0 = {[$:-1]};
		bins b1 = {[1:$]};
		option.weight = 1;
	 }

	//RS2 toggle bits
	rs2_val: coverpoint unsigned'(rv32m_trans.rs2_val) iff(rv32m_trans.trap==0) {
		wildcard bins b_1_0_0 	= (32'b???????????????????????????????1=>32'b???????????????????????????????0);
		wildcard bins b_1_0_1 	= (32'b??????????????????????????????1?=>32'b??????????????????????????????0?);
		wildcard bins b_1_0_2 	= (32'b?????????????????????????????1??=>32'b?????????????????????????????0??);
		wildcard bins b_1_0_3 	= (32'b????????????????????????????1???=>32'b????????????????????????????0???);
		wildcard bins b_1_0_4 	= (32'b???????????????????????????1????=>32'b???????????????????????????0????);
		wildcard bins b_1_0_5 	= (32'b??????????????????????????1?????=>32'b??????????????????????????0?????);
		wildcard bins b_1_0_6 	= (32'b?????????????????????????1??????=>32'b?????????????????????????0??????);
		wildcard bins b_1_0_7 	= (32'b????????????????????????1???????=>32'b????????????????????????0???????);
		wildcard bins b_1_0_8 	= (32'b???????????????????????1????????=>32'b???????????????????????0????????);
		wildcard bins b_1_0_9 	= (32'b??????????????????????1?????????=>32'b??????????????????????0?????????);
		wildcard bins b_1_0_10 	= (32'b?????????????????????1??????????=>32'b?????????????????????0??????????);
		wildcard bins b_1_0_11 	= (32'b????????????????????1???????????=>32'b????????????????????0???????????);
		wildcard bins b_1_0_12 	= (32'b???????????????????1????????????=>32'b???????????????????0????????????);
		wildcard bins b_1_0_13 	= (32'b??????????????????1?????????????=>32'b??????????????????0?????????????);
		wildcard bins b_1_0_14 	= (32'b?????????????????1??????????????=>32'b?????????????????0??????????????);
		wildcard bins b_1_0_15 	= (32'b????????????????1???????????????=>32'b????????????????0???????????????);
		wildcard bins b_1_0_16 	= (32'b???????????????1????????????????=>32'b???????????????0????????????????);
		wildcard bins b_1_0_17 	= (32'b??????????????1?????????????????=>32'b??????????????0?????????????????);
		wildcard bins b_1_0_18 	= (32'b?????????????1??????????????????=>32'b?????????????0??????????????????);
		wildcard bins b_1_0_19 	= (32'b????????????1???????????????????=>32'b????????????0???????????????????);
		wildcard bins b_1_0_20 	= (32'b???????????1????????????????????=>32'b???????????0????????????????????);
		wildcard bins b_1_0_21 	= (32'b??????????1?????????????????????=>32'b??????????0?????????????????????);
		wildcard bins b_1_0_22 	= (32'b?????????1??????????????????????=>32'b?????????0??????????????????????);
		wildcard bins b_1_0_23 	= (32'b????????1???????????????????????=>32'b????????0???????????????????????);
		wildcard bins b_1_0_24 	= (32'b???????1????????????????????????=>32'b???????0????????????????????????);
		wildcard bins b_1_0_25 	= (32'b??????1?????????????????????????=>32'b??????0?????????????????????????);
		wildcard bins b_1_0_26 	= (32'b?????1??????????????????????????=>32'b?????0??????????????????????????);
		wildcard bins b_1_0_27 	= (32'b????1???????????????????????????=>32'b????0???????????????????????????);
		wildcard bins b_1_0_28 	= (32'b???1????????????????????????????=>32'b???0????????????????????????????);
		wildcard bins b_1_0_29 	= (32'b??1?????????????????????????????=>32'b??0?????????????????????????????);
		wildcard bins b_1_0_30 	= (32'b?1??????????????????????????????=>32'b?0??????????????????????????????);
		wildcard bins b_1_0_31 	= (32'b1???????????????????????????????=>32'b0???????????????????????????????);
		wildcard bins b_0_1_0 	= (32'b???????????????????????????????0=>32'b???????????????????????????????1);
		wildcard bins b_0_1_1 	= (32'b??????????????????????????????0?=>32'b??????????????????????????????1?);
		wildcard bins b_0_1_2 	= (32'b?????????????????????????????0??=>32'b?????????????????????????????1??);
		wildcard bins b_0_1_3 	= (32'b????????????????????????????0???=>32'b????????????????????????????1???);
		wildcard bins b_0_1_4 	= (32'b???????????????????????????0????=>32'b???????????????????????????1????);
		wildcard bins b_0_1_5 	= (32'b??????????????????????????0?????=>32'b??????????????????????????1?????);
		wildcard bins b_0_1_6 	= (32'b?????????????????????????0??????=>32'b?????????????????????????1??????);
		wildcard bins b_0_1_7 	= (32'b????????????????????????0???????=>32'b????????????????????????1???????);
		wildcard bins b_0_1_8 	= (32'b???????????????????????0????????=>32'b???????????????????????1????????);
		wildcard bins b_0_1_9 	= (32'b??????????????????????0?????????=>32'b??????????????????????1?????????);
		wildcard bins b_0_1_10 	= (32'b?????????????????????0??????????=>32'b?????????????????????1??????????);
		wildcard bins b_0_1_11 	= (32'b????????????????????0???????????=>32'b????????????????????1???????????);
		wildcard bins b_0_1_12 	= (32'b???????????????????0????????????=>32'b???????????????????1????????????);
		wildcard bins b_0_1_13 	= (32'b??????????????????0?????????????=>32'b??????????????????1?????????????);
		wildcard bins b_0_1_14 	= (32'b?????????????????0??????????????=>32'b?????????????????1??????????????);
		wildcard bins b_0_1_15 	= (32'b????????????????0???????????????=>32'b????????????????1???????????????);
		wildcard bins b_0_1_16 	= (32'b???????????????0????????????????=>32'b???????????????1????????????????);
		wildcard bins b_0_1_17 	= (32'b??????????????0?????????????????=>32'b??????????????1?????????????????);
		wildcard bins b_0_1_18 	= (32'b?????????????0??????????????????=>32'b?????????????1??????????????????);
		wildcard bins b_0_1_19 	= (32'b????????????0???????????????????=>32'b????????????1???????????????????);
		wildcard bins b_0_1_20 	= (32'b???????????0????????????????????=>32'b???????????1????????????????????);
		wildcard bins b_0_1_21 	= (32'b??????????0?????????????????????=>32'b??????????1?????????????????????);
		wildcard bins b_0_1_22 	= (32'b?????????0??????????????????????=>32'b?????????1??????????????????????);
		wildcard bins b_0_1_23 	= (32'b????????0???????????????????????=>32'b????????1???????????????????????);
		wildcard bins b_0_1_24 	= (32'b???????0????????????????????????=>32'b???????1????????????????????????);
		wildcard bins b_0_1_25 	= (32'b??????0?????????????????????????=>32'b??????1?????????????????????????);
		wildcard bins b_0_1_26 	= (32'b?????0??????????????????????????=>32'b?????1??????????????????????????);
		wildcard bins b_0_1_27 	= (32'b????0???????????????????????????=>32'b????1???????????????????????????);
		wildcard bins b_0_1_28 	= (32'b???0????????????????????????????=>32'b???1????????????????????????????);
		wildcard bins b_0_1_29 	= (32'b??0?????????????????????????????=>32'b??1?????????????????????????????);
		wildcard bins b_0_1_30 	= (32'b?0??????????????????????????????=>32'b?1??????????????????????????????);
		wildcard bins b_0_1_31 	= (32'b0???????????????????????????????=>32'b1???????????????????????????????);
		option.weight = 1;
	 }

	//RS2 special values
	rs2_sp_val: coverpoint unsigned'(rv32m_trans.rs2_val) iff(rv32m_trans.trap==0) {
		bins b0 = {32'b0};
		bins b1 = {32'b00000000000000000000000000000001};
		bins b2 = {32'b11111111111111111111111111111111};
		bins b3 = {32'b01111111111111111111111111111111};
		bins b4 = {32'b10000000000000000000000000000000};
		bins b5 = {32'b10000000000000000000000000000001};
		option.weight = 1;
	 }

	//RS2 value sign
	rs2_val_sign: coverpoint rv32m_trans.rs2_val iff(rv32m_trans.trap==0) {
		bins b0 = {[$:-1]};
		bins b1 = {[1:$]};
		option.weight = 1;
	 }

	//war_hazard
	war_hazard_hit: coverpoint rv32m_trans.war_hazard_hit iff(rv32m_trans.trap==0) {
		bins b0 = {1};
		option.weight = 1;
	 }

	//waw_hazard
	waw_hazard_hit: coverpoint rv32m_trans.waw_hazard_hit iff(rv32m_trans.trap==0) {
		bins b0 = {1};
		option.weight = 1;
	 }

	//raw_hazard
	raw_hazard_hit: coverpoint rv32m_trans.raw_hazard_hit iff(rv32m_trans.trap==0) {
		bins b0 = {1};
		option.weight = 1;
	 }

	// base cross
	//MUL instruction crosspoints
	//Cross MUL instruction  and register assignment
	cr_mul_rs1_rs2_rd: cross mul,rs1_addr,rs2_addr,rd_addr {
		option.weight = 1;
	}

	//Cross MUL instruction  and RS1 toggle bits
	cr_mul_rs1_val: cross mul,rs1_val {
		option.weight = 1;
	}

	//Cross MUL instruction  and RS1 special values
	cr_mul_rs1_sp_val: cross mul,rs1_sp_val {
		option.weight = 1;
	}

	//Cross MUL instruction  and RS1 value sign
	cr_mul_rs1_val_sign: cross mul,rs1_val_sign {
		option.weight = 1;
	}

	//Cross MUL instruction  and RS2 toggle bits
	cr_mul_rs2_val: cross mul,rs2_val {
		option.weight = 1;
	}

	//Cross MUL instruction  and RS2 special values
	cr_mul_rs2_sp_val: cross mul,rs2_sp_val {
		option.weight = 1;
	}

	//Cross MUL instruction  and RS2 value sign
	cr_mul_rs2_val_sign: cross mul,rs2_val_sign {
		option.weight = 1;
	}

	//Cross MUL instruction  and RD toggle bits
	cr_mul_rd_val: cross mul,rd_val {
		option.weight = 1;
	}

	//Cross MUL instruction  and RD special values
	cr_mul_rd_sp_val: cross mul,rd_sp_val {
		option.weight = 1;
	}

	//Cross MUL instruction  and RD value sign
	cr_mul_rd_val_sign: cross mul,rd_val_sign {
		option.weight = 1;
	}

	//Cross MUL instruction  and WAR hazard
	cr_mul_war_hazard: cross mul,war_hazard_hit {
		option.weight = 1;
	}

	//Cross MUL instruction  and WAW hazard
	cr_mul_waw_hazard: cross mul,waw_hazard_hit {
		option.weight = 1;
	}

	//Cross MUL instruction  and RAW hazard
	cr_mul_raw_hazard: cross mul,raw_hazard_hit {
		option.weight = 1;
	}

	//MULH instruction crosspoints
	//Cross MULH instruction  and register assignment
	cr_mulh_rs1_rs2_rd: cross mulh,rs1_addr,rs2_addr,rd_addr {
		option.weight = 1;
	}

	//Cross MULH instruction  and RS1 toggle bits
	cr_mulh_rs1_val: cross mulh,rs1_val {
		option.weight = 1;
	}

	//Cross MULH instruction  and RS1 special values
	cr_mulh_rs1_sp_val: cross mulh,rs1_sp_val {
		option.weight = 1;
	}

	//Cross MULH instruction  and RS1 value sign
	cr_mulh_rs1_val_sign: cross mulh,rs1_val_sign {
		option.weight = 1;
	}

	//Cross MULH instruction  and RS2 toggle bits
	cr_mulh_rs2_val: cross mulh,rs2_val {
		option.weight = 1;
	}

	//Cross MULH instruction  and RS2 special values
	cr_mulh_rs2_sp_val: cross mulh,rs2_sp_val {
		option.weight = 1;
	}

	//Cross MULH instruction  and RS2 value sign
	cr_mulh_rs2_val_sign: cross mulh,rs2_val_sign {
		option.weight = 1;
	}

	//Cross MULH instruction  and RD toggle bits
	cr_mulh_rd_val: cross mulh,rd_val {
		option.weight = 1;
	}

	//Cross MULH instruction  and RD special values
	cr_mulh_rd_sp_val: cross mulh,rd_sp_val {
		option.weight = 1;
	}

	//Cross MULH instruction  and RD value sign
	cr_mulh_rd_val_sign: cross mulh,rd_val_sign {
		option.weight = 1;
	}

	//Cross MULH instruction  and WAR hazard
	cr_mulh_war_hazard: cross mulh,war_hazard_hit {
		option.weight = 1;
	}

	//Cross MULH instruction  and WAW hazard
	cr_mulh_waw_hazard: cross mulh,waw_hazard_hit {
		option.weight = 1;
	}

	//Cross MULH instruction  and RAW hazard
	cr_mulh_raw_hazard: cross mulh,raw_hazard_hit {
		option.weight = 1;
	}

	//MULHSU instruction crosspoints sign rs1,unsign rs2
	//Cross MULHSU instruction  and register assignment
	cr_mulhsu_rs1_rs2_rd: cross mulhsu,rs1_addr,rs2_addr,rd_addr {
		option.weight = 1;
	}

	//Cross MULHSU instruction  and RS1 toggle bits
	cr_mulhsu_rs1_val: cross mulhsu,rs1_val {
		option.weight = 1;
	}

	//Cross MULHSU instruction  and RS1 special values
	cr_mulhsu_rs1_sp_val: cross mulhsu,rs1_sp_val {
		option.weight = 1;
	}

	//Cross MULHSU instruction  and RS1 value sign
	cr_mulhsu_rs1_val_sign: cross mulhsu,rs1_val_sign {
		option.weight = 1;
	}

	//Cross MULHSU instruction  and RS2 toggle bits
	cr_mulhsu_rs2_val: cross mulhsu,rs2_val {
		option.weight = 1;
	}

	//Cross MULHSU instruction  and RS2 special values
	cr_mulhsu_rs2_sp_val: cross mulhsu,rs2_sp_val {
		option.weight = 1;
	}

	//Cross MULHSU instruction  and RD toggle bits
	cr_mulhsu_rd_val: cross mulhsu,rd_val {
		option.weight = 1;
	}

	//Cross MULHSU instruction  and RD special values
	cr_mulhsu_rd_sp_val: cross mulhsu,rd_sp_val {
		option.weight = 1;
	}

	//Cross MULHSU instruction  and RD value sign
	cr_mulhsu_rd_val_sign: cross mulhsu,rd_val_sign {
		option.weight = 1;
	}

	//Cross MULHSU instruction  and WAR hazard
	cr_mulhsu_war_hazard: cross mulhsu,war_hazard_hit {
		option.weight = 1;
	}

	//Cross MULHSU instruction  and WAW hazard
	cr_mulhsu_waw_hazard: cross mulhsu,waw_hazard_hit {
		option.weight = 1;
	}

	//Cross MULHSU instruction  and RAW hazard
	cr_mulhsu_raw_hazard: cross mulhsu,raw_hazard_hit {
		option.weight = 1;
	}

	//MULHU instruction  unsign
	//Cross MULHU instruction  and register assignment
	cr_mulhu_rs1_rs2_rd: cross mulhu,rs1_addr,rs2_addr,rd_addr {
		option.weight = 1;
	}

	//Cross MULHU instruction  and RS1 toggle bits
	cr_mulhu_rs1_val: cross mulhu,rs1_val {
		option.weight = 1;
	}

	//Cross MULHU instruction  and RS1 special values
	cr_mulhu_rs1_sp_val: cross mulhu,rs1_sp_val {
		option.weight = 1;
	}

	//Cross MULHU instruction  and RS2 toggle bits
	cr_mulhu_rs2_val: cross mulhu,rs2_val {
		option.weight = 1;
	}

	//Cross MULHU instruction  and RS2 special values
	cr_mulhu_rs2_sp_val: cross mulhu,rs2_sp_val {
		option.weight = 1;
	}

	//Cross MULHU instruction  and RD toggle bits
	cr_mulhu_rd_val: cross mulhu,rd_val {
		option.weight = 1;
	}

	//Cross MULHU instruction  and RD special values
	cr_mulhu_rd_sp_val: cross mulhu,rd_sp_val {
		option.weight = 1;
	}

	//Cross MULHU instruction  and WAR hazard
	cr_mulhu_war_hazard: cross mulhu,war_hazard_hit {
		option.weight = 1;
	}

	//Cross MULHU instruction  and WAW hazard
	cr_mulhu_waw_hazard: cross mulhu,waw_hazard_hit {
		option.weight = 1;
	}

	//Cross MULHU instruction  and RAW hazard
	cr_mulhu_raw_hazard: cross mulhu,raw_hazard_hit {
		option.weight = 1;
	}

	//DIV instruction crosspoints
	//Cross DIV instruction  and register assignment
	cr_div_rs1_rs2_rd: cross div,rs1_addr,rs2_addr,rd_addr {
		option.weight = 1;
	}

	//Cross DIV instruction  and RS1 toggle bits
	cr_div_rs1_val: cross div,rs1_val {
		option.weight = 1;
	}

	//Cross DIV instruction  and RS1 special values
	cr_div_rs1_sp_val: cross div,rs1_sp_val {
		option.weight = 1;
	}

	//Cross DIV instruction  and RS1 value sign
	cr_div_rs1_val_sign: cross div,rs1_val_sign {
		option.weight = 1;
	}

	//Cross DIV instruction  and RS2 toggle bits
	cr_div_rs2_val: cross div,rs2_val {
		option.weight = 1;
	}

	//Cross DIV instruction  and RS2 special values
	cr_div_rs2_sp_val: cross div,rs2_sp_val {
		option.weight = 1;
	}

	//Cross DIV instruction  and RS2 value sign
	cr_div_rs2_val_sign: cross div,rs2_val_sign {
		option.weight = 1;
	}

	//Cross DIV instruction  and RD toggle bits
	cr_div_rd_val: cross div,rd_val {
		option.weight = 1;
	}

	//Cross DIV instruction  and RD special values
	cr_div_rd_sp_val: cross div,rd_sp_val {
		option.weight = 1;
	}

	//Cross DIV instruction  and RD value sign
	cr_div_rd_val_sign: cross div,rd_val_sign {
		option.weight = 1;
	}

	//Cross DIV instruction  and WAR hazard
	cr_div_war_hazard: cross div,war_hazard_hit {
		option.weight = 1;
	}

	//Cross DIV instruction  and WAW hazard
	cr_div_waw_hazard: cross div,waw_hazard_hit {
		option.weight = 1;
	}

	//Cross DIV instruction  and RAW hazard
	cr_div_raw_hazard: cross div,raw_hazard_hit {
		option.weight = 1;
	}

	//overflow -2^31 / -1
	cr_div_overflow: cross div,rs1_sp_val,rs2_sp_val {
		option.weight = 1;
	}

	//x / 0 = -1
	cr_div_division_by_zero: cross div,rd_sp_val,rs2_sp_val {
		bins div_zero = binsof(div) intersect {DIV} && binsof(rd_sp_val) intersect {32'b11111111111111111111111111111111} && binsof(rs2_sp_val) intersect{32'b0};
		option.weight = 1;
	}
	//DIVU instruction  unsign
	//Cross DIVU instruction  and register assignment
	cr_divu_rs1_rs2_rd: cross divu,rs1_addr,rs2_addr,rd_addr {
		option.weight = 1;
	}

	//Cross DIVU instruction  and RS1 toggle bits
	cr_divu_rs1_val: cross divu,rs1_val {
		option.weight = 1;
	}

	//Cross DIVU instruction  and RS1 special values
	cr_divu_rs1_sp_val: cross divu,rs1_sp_val {
		option.weight = 1;
	}

	//Cross DIVU instruction  and RS2 toggle bits
	cr_divu_rs2_val: cross divu,rs2_val {
		option.weight = 1;
	}

	//Cross DIVU instruction  and RS2 special values
	cr_divu_rs2_sp_val: cross divu,rs2_sp_val {
		option.weight = 1;
	}

	//Cross DIVU instruction  and RD toggle bits
	cr_divu_rd_val: cross divu,rd_val {
		option.weight = 1;
	}

	//Cross DIVU instruction  and RD special values
	cr_divu_rd_sp_val: cross divu,rd_sp_val {
		option.weight = 1;
	}

	//Cross DIVU instruction  and WAR hazard
	cr_divu_war_hazard: cross divu,war_hazard_hit {
		option.weight = 1;
	}

	//Cross DIVU instruction  and WAW hazard
	cr_divu_waw_hazard: cross divu,waw_hazard_hit {
		option.weight = 1;
	}

	//Cross DIVU instruction  and RAW hazard
	cr_divu_raw_hazard: cross divu,raw_hazard_hit {
		option.weight = 1;
	}

	//x / 0 = -1
	cr_divu_division_by_zero: cross divu,rd_sp_val,rs2_sp_val {
		bins divu_zero = binsof(divu) intersect {DIVU} && binsof(rd_sp_val) intersect {32'b11111111111111111111111111111111} && binsof(rs2_sp_val) intersect{32'b0};
		option.weight = 1;
	}
	//REM instruction crosspoints
	//Cross REM instruction  and register assignment
	cr_rem_rs1_rs2_rd: cross rem,rs1_addr,rs2_addr,rd_addr {
		option.weight = 1;
	}

	//Cross REM instruction  and RS1 toggle bits
	cr_rem_rs1_val: cross rem,rs1_val {
		option.weight = 1;
	}

	//Cross REM instruction  and RS1 special values
	cr_rem_rs1_sp_val: cross rem,rs1_sp_val {
		option.weight = 1;
	}

	//Cross REM instruction  and RS1 value sign
	cr_rem_rs1_val_sign: cross rem,rs1_val_sign {
		option.weight = 1;
	}

	//Cross REM instruction  and RS2 toggle bits
	cr_rem_rs2_val: cross rem,rs2_val {
		option.weight = 1;
	}

	//Cross REM instruction  and RS2 special values
	cr_rem_rs2_sp_val: cross rem,rs2_sp_val {
		option.weight = 1;
	}

	//Cross REM instruction  and RS2 value sign
	cr_rem_rs2_val_sign: cross rem,rs2_val_sign {
		option.weight = 1;
	}

	//Cross REM instruction  and RD toggle bits
	cr_rem_rd_val: cross rem,rd_val {
		option.weight = 1;
	}

	//Cross REM instruction  and RD special values
	cr_rem_rd_sp_val: cross rem,rd_sp_val {
		option.weight = 1;
	}

	//Cross REM instruction  and RD value sign
	cr_rem_rd_val_sign: cross rem,rd_val_sign {
		option.weight = 1;
	}

	//Cross REM instruction  and WAR hazard
	cr_rem_war_hazard: cross rem,war_hazard_hit {
		option.weight = 1;
	}

	//Cross REM instruction  and WAW hazard
	cr_rem_waw_hazard: cross rem,waw_hazard_hit {
		option.weight = 1;
	}

	//Cross REM instruction  and RAW hazard
	cr_rem_raw_hazard: cross rem,raw_hazard_hit {
		option.weight = 1;
	}

	//x % 0 = x
	cr_rem_division_by_zero: cross rem,rs2_sp_val {
		bins rem_zero = binsof(rem) intersect {REM}&& binsof(rs2_sp_val) intersect{32'b0};
		option.weight = 1;
	}
	//REMU instruction  unsign
	//Cross REMU instruction  and register assignment
	cr_remu_rs1_rs2_rd: cross remu,rs1_addr,rs2_addr,rd_addr {
		option.weight = 1;
	}

	//Cross REMU instruction  and RS1 toggle bits
	cr_remu_rs1_val: cross remu,rs1_val {
		option.weight = 1;
	}

	//Cross REMU instruction  and RS1 special values
	cr_remu_rs1_sp_val: cross remu,rs1_sp_val {
		option.weight = 1;
	}

	//Cross REMU instruction  and RS2 toggle bits
	cr_remu_rs2_val: cross remu,rs2_val {
		option.weight = 1;
	}

	//Cross REMU instruction  and RS2 special values
	cr_remu_rs2_sp_val: cross remu,rs2_sp_val {
		option.weight = 1;
	}

	//Cross REMU instruction  and RD toggle bits
	cr_remu_rd_val: cross remu,rd_val {
		option.weight = 1;
	}

	//Cross REMU instruction  and RD special values
	cr_remu_rd_sp_val: cross remu,rd_sp_val {
		option.weight = 1;
	}

	//Cross REMU instruction  and WAR hazard
	cr_remu_war_hazard: cross remu,war_hazard_hit {
		option.weight = 1;
	}

	//Cross REMU instruction  and WAW hazard
	cr_remu_waw_hazard: cross remu,waw_hazard_hit {
		option.weight = 1;
	}

	//Cross REMU instruction  and RAW hazard
	cr_remu_raw_hazard: cross remu,raw_hazard_hit {
		option.weight = 1;
	}

	//x % 0 = x
	cr_remu_division_by_zero: cross remu,rs2_sp_val {
		bins remu_zero = binsof(remu) intersect {REMU}&& binsof(rs2_sp_val) intersect{32'b0};
		option.weight = 1;
	}

endgroup
